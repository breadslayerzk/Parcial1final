library verilog;
use verilog.vl_types.all;
entity peaje_electronico_vlg_vec_tst is
end peaje_electronico_vlg_vec_tst;
